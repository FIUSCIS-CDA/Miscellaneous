///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: Miscellaneous
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"


//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing Decoder_32
reg[4:0] A;
wire[31:0] Q;
Decoder_32 myDecoder(
        .A(A),
        .Q0(Q[0]),.Q1(Q[1]),.Q2(Q[2]),.Q3(Q[3]),.Q4(Q[4]),.Q5(Q[5]),.Q6(Q[6]),.Q7(Q[7]),
        .Q8(Q[8]),.Q9(Q[9]),.Q10(Q[10]),.Q11(Q[11]),.Q12(Q[12]),.Q13(Q[13]),.Q14(Q[14]),.Q15(Q[15]),
        .Q16(Q[16]),.Q17(Q[17]),.Q18(Q[18]),.Q19(Q[19]),.Q20(Q[20]),.Q21(Q[21]),.Q22(Q[22]),.Q23(Q[23]),
        .Q24(Q[24]),.Q25(Q[25]),.Q26(Q[26]),.Q27(Q[27]),.Q28(Q[28]),.Q29(Q[29]),.Q30(Q[30]),.Q31(Q[31])
);

//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing Encoder_32
reg[31:0] AENC;
wire[4:0] QENC;
Encoder_32 myEncoder(
        .A0(AENC[0]),.A1(AENC[1]),.A2(AENC[2]),.A3(AENC[3]),.A4(AENC[4]),.A5(AENC[5]),.A6(AENC[6]),.A7(AENC[7]),
        .A8(AENC[8]),.A9(AENC[9]),.A10(AENC[10]),.A11(AENC[11]),.A12(AENC[12]),.A13(AENC[13]),.A14(AENC[14]),.A15(AENC[15]),
        .A16(AENC[16]),.A17(AENC[17]),.A18(AENC[18]),.A19(AENC[19]),.A20(AENC[20]),.A21(AENC[21]),.A22(AENC[22]),.A23(AENC[23]),
        .A24(AENC[24]),.A25(AENC[25]),.A26(AENC[26]),.A27(AENC[27]),.A28(AENC[28]),.A29(AENC[29]),.A30(AENC[30]),.A31(AENC[31]),
        .Q(QENC));
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing SameBit
reg Ain;
wire Aout;
SameBit mySame(.Ain(Ain), .Aout(Aout));
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing SPLICE_PCJ
reg[25:0] ir25_0;
reg[3:0] pc31_28;
wire[31:0] Y; 
SPLICE_PCJ mySplicer(.ir25_0(ir25_0), .pc31_28(pc31_28), .Y(Y));
//////////////////////////////////////////////////////////////////////////////////////////////////////

initial begin 
////////////////////////////////////////////////////////////////////////////////////////
// 

A = 5'b01101;
AENC = 32'b00000010000000000000000000000000;
Ain=0;
pc31_28=4'b0110; ir25_0=26'b00001100011000000001101011;  
#10;
   $display("Testing: A=%b", A);
verifyEqual32(Q, 2**A);
   $display("Testing: AENC=%b", AENC);
verifyEqual5(QENC, 25);
$display("Testing: Ain=0");
verifyEqual(Aout, Ain);
$display("Test: pc31_28=0110, ir25_0=b00001100011000000001101011");
verifyEqual32(Y, {pc31_28, ir25_0, 2'b00});


// Encoder_32

////////////////////////////////////////////////////////////////////////////////////////
 
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule